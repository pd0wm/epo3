configuration sr_demux8_inv_sr_demux8_inv_behav_cfg of sr_demux8_inv is
   for sr_demux8_inv_behav
   end for;
end sr_demux8_inv_sr_demux8_inv_behav_cfg;


