configuration vga_demux_vga_demux_behav_cfg of vga_demux is
   for vga_demux_behav
   end for;
end vga_demux_vga_demux_behav_cfg;


