configuration bit4_bit4_behav_cfg of bit4 is
   for bit4_behav
   end for;
end bit4_bit4_behav_cfg;


