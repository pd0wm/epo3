configuration cs_tri7_cs_tri7_behav_cfg of cs_tri7 is
   for cs_tri7_behav
   end for;
end cs_tri7_cs_tri7_behav_cfg;


