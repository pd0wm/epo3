configuration controller_calc_controller_calc_arch_cfg of controller_calc is
   for controller_calc_arch
   end for;
end controller_calc_controller_calc_arch_cfg;


