configuration piece_lut_extracted_cfg of piece_lut is
   for extracted
   end for;
end piece_lut_extracted_cfg;


