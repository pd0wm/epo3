configuration debounce_behaviour_cfg of debounce is
   for behaviour
   end for;
end debounce_behaviour_cfg;


