configuration top_level2_tb_top_level2_tb_arch_cfg of top_level2_tb is
   for top_level2_tb_arch
      for all: top_level2 use configuration work.top_level2_top_level2_struc_cfg;
      end for;
   end for;
end top_level2_tb_top_level2_tb_arch_cfg;


