configuration de_piece_behaviour_cfg of de_piece is
   for behaviour
   end for;
end de_piece_behaviour_cfg;


