configuration rom_tb_behaviour_cfg of rom_tb is
   for rom_tb_behaviour
      for all: rom use configuration work.rom_behaviour_cfg;
      end for;
   end for;
end rom_tb_behaviour_cfg;


