configuration vga_counter_10bit_vga_counter_10bit_behav_cfg of vga_counter_10bit is
   for vga_counter_10bit_behav
   end for;
end vga_counter_10bit_vga_counter_10bit_behav_cfg;


