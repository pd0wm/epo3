configuration timer_behaviour_cfg of timer is
   for behaviour
   end for;
end timer_behaviour_cfg;


