configuration timer_synthesised_cfg of timer is
   for synthesised
   end for;
end timer_synthesised_cfg;


