configuration vga_trans_reset_vga_trans_reset_arch_cfg of vga_trans_reset is
   for vga_trans_reset_arch
   end for;
end vga_trans_reset_vga_trans_reset_arch_cfg;


