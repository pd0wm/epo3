library IEEE;
use IEEE.std_logic_1164.ALL;

entity top_level_tb is
end top_level_tb;
