configuration sr_tower_tb_sr_tower_tb_behav_cfg of sr_tower_tb is
   for sr_tower_tb_behav
      for all: sr_tower use configuration work.sr_tower_sr_tower_behav_cfg;
      end for;
   end for;
end sr_tower_tb_sr_tower_tb_behav_cfg;


