configuration vga_score_trans_vga_score_trans_arch_cfg of vga_score_trans is
   for vga_score_trans_arch
      for all: vga_counter_3bit use configuration work.vga_counter_3bit_vga_counter_3bit_behav_cfg;
      end for;
   end for;
end vga_score_trans_vga_score_trans_arch_cfg;


