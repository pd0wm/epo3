library ieee;
use ieee.std_logic_1164.all;
entity controller_calc is
	port(
		clk               : in  std_logic;
		rst               : in  std_logic

	);
end controller_calc;



