configuration extracted of sr_if_tb is
   for sr_if_tb_behav
      for all: sr_if use configuration work.sr_if_extracted_cfg;
      end for;
   end for;
end extracted;


