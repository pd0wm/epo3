configuration check_mask_synthesised_cfg of check_mask is
   for synthesised
   end for;
end check_mask_synthesised_cfg;


