configuration tri_buff_synthesised_cfg of tri_buff is
   for synthesised
   end for;
end tri_buff_synthesised_cfg;


