configuration vga_np_trans_vga_np_trans_arch_cfg of vga_np_trans is
   for vga_np_trans_arch
      for all: vga_counter_8bitset use configuration work.vga_counter_8bitset_vga_counter_8bitset_behav_cfg;
      end for;
   end for;
end vga_np_trans_vga_np_trans_arch_cfg;


