configuration vga_score_trans_vga_score_trans_arch_cfg of vga_score_trans is
   for vga_score_trans_arch
   end for;
end vga_score_trans_vga_score_trans_arch_cfg;


