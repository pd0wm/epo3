configuration rom_mux2_behaviour_cfg of rom_mux2 is
   for rom_mux2_behaviour
   end for;
end rom_mux2_behaviour_cfg;


