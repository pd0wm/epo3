configuration score_behaviour_cfg of score is
   for behaviour
   end for;
end score_behaviour_cfg;


