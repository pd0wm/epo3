configuration draw_score_synthesised_cfg of draw_score is
   for synthesised
   end for;
end draw_score_synthesised_cfg;


