configuration vga_np_check_vga_np_check_arch_cfg of vga_np_check is
   for vga_np_check_arch
   end for;
end vga_np_check_vga_np_check_arch_cfg;


