configuration piece_lut_synthesised_cfg of piece_lut is
   for synthesised
   end for;
end piece_lut_synthesised_cfg;


