configuration vga_counter_vga_counter_behav_cfg of vga_counter is
   for vga_counter_behav
   end for;
end vga_counter_vga_counter_behav_cfg;


