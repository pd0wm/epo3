configuration checkmask_tb_behaviour_ext_fg of checkmask_tb is
   for checkmask_tb_behaviour
      for all: checkmask use configuration work.checkmask_extracted_cfg;
      end for;
   end for;
end checkmask_tb_behaviour_ext_fg;


