


library ieee;
use ieee.std_logic_1164.all;

package vga_params2 is

	
end vga_params2;

package body vga_params2 is
end vga_params2;






