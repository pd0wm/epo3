configuration checkmask_extracted_cfg of checkmask is
   for extracted
   end for;
end checkmask_extracted_cfg;


