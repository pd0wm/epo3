library IEEE;
use IEEE.std_logic_1164.ALL;

entity clearshift_tb is
end clearshift_tb;


