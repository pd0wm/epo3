library ieee;
use ieee.std_logic_1164.all;

entity cs_defset2 is
	port(
		en   : in  std_logic;
		out1 : out std_logic;
		out2 : out std_logic
	);
end entity;