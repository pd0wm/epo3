library IEEE;
use IEEE.std_logic_1164.ALL;

architecture fake_ram_arch of fake_ram is
begin
end fake_ram_arch;


