configuration vga_np_trans_reset_vga_np_trans_reset_arch_cfg of vga_np_trans_reset is
   for vga_np_trans_reset_arch
      for all: vga_counter_2bit use configuration work.vga_counter_2bit_vga_counter_2bit_behav_cfg;
      end for;
   end for;
end vga_np_trans_reset_vga_np_trans_reset_arch_cfg;


