configuration bit4_tb_bit4_tb_behav_cfg of bit4_tb is
   for bit4_tb_behav
      for all: bit4 use configuration work.bit4_bit4_behav_cfg;
      end for;
   end for;
end bit4_tb_bit4_tb_behav_cfg;


