configuration vga_field_trans_reset_vga_field_trans_reset_arch_cfg of vga_field_trans_reset is
   for vga_field_trans_reset_arch
      for all: vga_counter_4bit use configuration work.vga_counter_4bit_vga_counter_4bit_behav_cfg;
      end for;
   end for;
end vga_field_trans_reset_vga_field_trans_reset_arch_cfg;


