configuration vga_counter_5bit_vga_counter_5bit_behav_cfg of vga_counter_5bit is
   for vga_counter_5bit_behav
   end for;
end vga_counter_5bit_vga_counter_5bit_behav_cfg;


