configuration sr_demux4_inv_sr_demux4_inv_behav_cfg of sr_demux4_inv is
   for sr_demux4_inv_behav
   end for;
end sr_demux4_inv_sr_demux4_inv_behav_cfg;


