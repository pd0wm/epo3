configuration score_extracted_cfg of score is
   for extracted
   end for;
end score_extracted_cfg;


