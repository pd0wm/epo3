configuration cs_compare_tb_old_cs_compare_tb_behav_cfg of cs_compare_tb_old is
   for cs_compare_tb_behav


