configuration score_synthesised_cfg of score is
   for synthesised
   end for;
end score_synthesised_cfg;


