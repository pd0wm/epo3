library IEEE;
use IEEE.std_logic_1164.ALL;

entity rom_tb is
end rom_tb;


