configuration controller_controller_arch_cfg of controller is
   for controller_arch
   end for;
end controller_controller_arch_cfg;


