library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.vga_params.all;

entity vga_tb is
	constant clk_period : time := 20 ns;
end entity;

architecture vga_tb_arch of vga_tb is
	component vga
		port(clk      : in  std_logic;
			 rst      : in  std_logic;
			 mem_addr : out std_logic_vector(mem_addr_len - 1 downto 0);
			 data     : in  std_logic;
			 h_sync   : out std_logic;
			 v_sync   : out std_logic;
			 red      : out std_logic;
			 green    : out std_logic;
			 blue     : out std_logic);
	end component vga;

	signal clk, rst, data : std_logic;
	signal h_sync, v_sync : std_logic;
	signal ram_addr       : std_logic_vector(6 downto 0);

	signal r, g, b : std_logic;

begin
	uut : vga
		port map(clk      => clk,
			     rst      => rst,
			     mem_addr => ram_addr,
			     data     => data,
			     h_sync   => h_sync,
			     v_sync   => v_sync,
			     red      => r,
			     green    => g,
			     blue     => b);
	clock : process
	begin
		clk <= '1';
		wait for clk_period / 2;
		clk <= '0';
		wait for clk_period / 2;
	end process;

	data_lut : process(clk, rst)
		variable addr : integer;
	begin
		if (rst = '1') then
			data <= '0';
		elsif (clk'event and clk = '1') then
			addr := to_integer(unsigned(ram_addr));
			data <= '0';

			if (
				addr = 5 or addr = 6 or addr = 9 or addr = 10
			) then
				data <= '1';
			end if;
		end if;
	end process;

	rst <= '1', '0' after clk_period;
end;



