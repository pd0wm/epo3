configuration vga_sync_vga_sync_arch_cfg of vga_sync is
   for vga_sync_arch
   end for;
end vga_sync_vga_sync_arch_cfg;


