configuration sr_demux5_sr_demux5_behav_cfg of sr_demux5 is
   for sr_demux5_behav
   end for;
end sr_demux5_sr_demux5_behav_cfg;


