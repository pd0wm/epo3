configuration timer_extracted_cfg of timer is
   for extracted
   end for;
end timer_extracted_cfg;


