library IEEE;
use IEEE.std_logic_1164.ALL;

entity ram_simple is
end ram_simple;


