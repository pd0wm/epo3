library IEEE;
use IEEE.std_logic_1164.ALL;

entity piece_lut_tb is
end piece_lut_tb;


