configuration clearandshift_extracted_cfg of clearandshift is
   for extracted
   end for;
end clearandshift_extracted_cfg;


