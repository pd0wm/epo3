configuration cs_adder7_cs_addr7_behav_cfg of cs_adder7 is
   for cs_addr7_behav
   end for;
end cs_adder7_cs_addr7_behav_cfg;


