configuration log_behaviour_cfg of log is
   for behaviour
   end for;
end log_behaviour_cfg;


