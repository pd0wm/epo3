configuration vga_field_trans_vga_field_trans_arch_cfg of vga_field_trans is
   for vga_field_trans_arch
   end for;
end vga_field_trans_vga_field_trans_arch_cfg;


