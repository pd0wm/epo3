configuration vga_score_check_vga_score_check_arch_cfg of vga_score_check is
   for vga_score_check_arch
   end for;
end vga_score_check_vga_score_check_arch_cfg;


