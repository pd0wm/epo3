configuration cs_defset2_cs_defset2_behav_cfg of cs_defset2 is
   for cs_defset2_behav
   end for;
end cs_defset2_cs_defset2_behav_cfg;


