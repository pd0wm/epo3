configuration cs_shift_extracted_cfg of cs_shift is
   for extracted
   end for;
end cs_shift_extracted_cfg;


