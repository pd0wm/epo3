configuration check_mask_behaviour_cfg of check_mask is
   for check_mask_behaviour
   end for;
end check_mask_behaviour_cfg;


