configuration top_top_level_tb_behaviour_cfg of top_top_level_tb is
   for behaviour
      for all: top_top_level use configuration work.top_top_level_top_top_level_struc_cfg;
      end for;
   end for;
end top_top_level_tb_behaviour_cfg;


