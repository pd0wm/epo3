configuration demux5_demux5_behav_cfg of demux5 is
   for demux5_behav
   end for;
end demux5_demux5_behav_cfg;


