configuration cs_7bc_cs_7bc_arch_cfg of cs_7bc is
   for cs_7bc_arch
   end for;
end cs_7bc_cs_7bc_arch_cfg;


