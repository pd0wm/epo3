library IEEE;
use IEEE.std_logic_1164.ALL;

entity fake_ram is
end fake_ram;


