configuration checkmask_behaviour_cfg of checkmask is
   for checkmask_behaviour
   end for;
end checkmask_behaviour_cfg;


