configuration vga_np_trans_reset_vga_np_trans_reset_arch_cfg of vga_np_trans_reset is
   for vga_np_trans_reset_arch
   end for;
end vga_np_trans_reset_vga_np_trans_reset_arch_cfg;


