configuration dec8_dec8_behav_cfg of dec8 is
   for dec8_behav
   end for;
end dec8_dec8_behav_cfg;


