library ieee;
use ieee.std_logic_1164.all;

package typedef is
	type mem is array (0 to 2**8-1) of std_logic;
end typedef;

package body typedef is
end typedef;