configuration vga_triggers_vga_triggers_arch_cfg of vga_triggers is
   for vga_triggers_arch
   end for;
end vga_triggers_vga_triggers_arch_cfg;


