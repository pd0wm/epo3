configuration vga_counter_resets_vga_counter_resets_behav_cfg of vga_counter_resets is
   for vga_counter_resets_behav
   end for;
end vga_counter_resets_vga_counter_resets_behav_cfg;


