library ieee;
use ieee.std_logic_1164.all;

entity ram_simple is
	port(
		clk             : in    std_logic;
		rst             : in    std_logic;

		rw_addr         : in    std_logic_vector(7 downto 0);
		rw_data         : inout std_logic;
		rw_write_enable : in    std_logic;

		ro_addr         : in    std_logic_vector(7 downto 0);
		ro_out          : out   std_logic
	);

end ram_simple;

