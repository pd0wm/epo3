library ieee;
use ieee.std_logic_1164.all;

package mem is
	type mem is array (0 to 2**5-1) of std_logic;
end mem;

package body mem is
end mem;