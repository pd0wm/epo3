configuration log_synthesised_cfg of log is
   for synthesised
   end for;
end log_synthesised_cfg;


