library IEEE;
use IEEE.std_logic_1164.ALL;

entity score_tb is
end score_tb;


