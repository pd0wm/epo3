library IEEE;
use IEEE.std_logic_1164.ALL;

architecture depiece_simple_arch of depiece_simple is
begin
end depiece_simple_arch;


