configuration log_score_tb_behaviour_cfg of log_score_tb is
   for behaviour
      for all: log_score use configuration work.log_score_behaviour_cfg;
      end for;
   end for;
end log_score_tb_behaviour_cfg;


