configuration check_mask_extracted_cfg of check_mask is
   for extracted
   end for;
end check_mask_extracted_cfg;


