configuration npg_ff_behaviour_cfg of npg_ff is
   for behaviour
   end for;
end npg_ff_behaviour_cfg;


