configuration timer_det_timer_det_arch_cfg of timer_det is
   for timer_det_arch
   end for;
end timer_det_timer_det_arch_cfg;


