configuration cs_7bcws_cs_7bcws_behav_cfg of cs_7bcws is
   for cs_7bcws_behav
   end for;
end cs_7bcws_cs_7bcws_behav_cfg;


