configuration vga_tb_vga_tb_arch_cfg of vga_tb is
   for vga_tb_arch
   end for;
end vga_tb_vga_tb_arch_cfg;


