configuration adder_y_behaviour_cfg of adder_y is
   for behaviour
   end for;
end adder_y_behaviour_cfg;


