configuration vga_trans_vga_trans_arch_cfg of vga_trans is
   for vga_trans_arch
   end for;
end vga_trans_vga_trans_arch_cfg;


