configuration clearandshift_behaviour_cfg of clearandshift is
   for clearandshift_behaviour
   end for;
end clearandshift_behaviour_cfg;


