configuration vga_field_trans_reset_vga_field_trans_reset_arch_cfg of vga_field_trans_reset is
   for vga_field_trans_reset_arch
   end for;
end vga_field_trans_reset_vga_field_trans_reset_arch_cfg;


