configuration sr_bit4_sr_bit4_behav_cfg of sr_bit4 is
   for sr_bit4_behav
   end for;
end sr_bit4_sr_bit4_behav_cfg;


