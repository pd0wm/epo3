configuration log_score_extracted_cfg of log_score is
   for extracted
   end for;
end log_score_extracted_cfg;


