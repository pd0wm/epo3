configuration sr_if_extracted_cfg of sr_if is
   for extracted
   end for;
end sr_if_extracted_cfg;


