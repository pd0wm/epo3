library IEEE;
use IEEE.std_logic_1164.ALL;

architecture controller_arch of controller is
begin
end controller_arch;


