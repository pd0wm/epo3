configuration ram_simple_ram_simple_arch_cfg of ram_simple is
   for ram_simple_arch
   end for;
end ram_simple_ram_simple_arch_cfg;


