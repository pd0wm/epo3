library IEEE;
use IEEE.std_logic_1164.ALL;

architecture ram_simple_arch of ram_simple is
begin
end ram_simple_arch;


