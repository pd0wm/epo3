configuration vga_read_vga_read_behav_cfg of vga_read is
   for vga_read_behav
   end for;
end vga_read_vga_read_behav_cfg;


