configuration vga_np_trans_vga_np_trans_arch_cfg of vga_np_trans is
   for vga_np_trans_arch
   end for;
end vga_np_trans_vga_np_trans_arch_cfg;


