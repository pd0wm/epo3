library IEEE;
use IEEE.std_logic_1164.ALL;

entity timer_tb is
end timer_tb;


