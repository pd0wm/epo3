library IEEE;
use IEEE.std_logic_1164.ALL;

entity npg_tb is
end npg_tb;


