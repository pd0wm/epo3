configuration ram_fix_ram_fix_behav_cfg of ram_fix is
   for ram_fix_behav
   end for;
end ram_fix_ram_fix_behav_cfg;


