configuration vga_extracted_cfg of vga is
   for extracted
   end for;
end vga_extracted_cfg;


