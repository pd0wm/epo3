configuration tri_buff_behaviour_cfg of tri_buff is
   for behaviour
   end for;
end tri_buff_behaviour_cfg;


