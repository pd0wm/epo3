configuration vga_counter_4bit_vga_counter_4bit_behav_cfg of vga_counter_4bit is
   for vga_counter_4bit_behav
   end for;
end vga_counter_4bit_vga_counter_4bit_behav_cfg;


