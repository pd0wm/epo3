library IEEE;
use IEEE.std_logic_1164.ALL;

entity de_piece_tb is
end de_piece_tb;


