configuration controller_tb_behaviour_cfg of controller_tb is
   for behaviour
      for all: controller use configuration work.controller_controller_arch_cfg;
      end for;
   end for;
end controller_tb_behaviour_cfg;


