configuration adder_x_behaviour_cfg of adder_x is
   for behaviour
   end for;
end adder_x_behaviour_cfg;


