configuration de_piece_testbench_behaviour_cfg of de_piece_testbench is
   for behaviour
      for all: de_piece use configuration work.de_piece_behaviour_cfg;
      end for;
   end for;
end de_piece_testbench_behaviour_cfg;


