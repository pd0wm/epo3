configuration cs_compare_comb_cs_compare_comb_behav_cfg of cs_compare_comb is
   for cs_compare_comb_behav
   end for;
end cs_compare_comb_cs_compare_comb_behav_cfg;


