configuration demux8_inv_demux8_inv_behav_cfg of demux8_inv is
   for demux8_inv_behav
   end for;
end demux8_inv_demux8_inv_behav_cfg;


