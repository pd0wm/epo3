configuration sr_dec8_sr_dec8_behav_cfg of sr_dec8 is
   for sr_dec8_behav
   end for;
end sr_dec8_sr_dec8_behav_cfg;


