configuration sr_mux5_sr_mux5_behav_cfg of sr_mux5 is
   for sr_mux5_behav
   end for;
end sr_mux5_sr_mux5_behav_cfg;


