configuration log_score_syn_tb_behaviour_cfg of log_score_tb is
   for behaviour
      for all: log_score use configuration work.log_score_synthesised_cfg;
      end for;
   end for;
end log_score_syn_tb_behaviour_cfg;


