configuration piece_lut_tb_behaviour_syn_cfg of piece_lut_tb is
   for piece_lut_tb_behaviour
      for all: piece_lut use configuration work.piece_lut_behaviour_cfg;
      end for;
   end for;
end piece_lut_tb_behaviour_syn_cfg;


