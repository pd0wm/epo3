configuration top_top_level_top_top_level_struc_cfg of top_top_level is
   for top_top_level_struc
      for all: top_level2 use configuration work.top_level2_top_level2_struc_cfg;
      end for;
   end for;
end top_top_level_top_top_level_struc_cfg;


