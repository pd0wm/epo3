configuration checkmask_synthesised_cfg of checkmask is
   for synthesised
   end for;
end checkmask_synthesised_cfg;


