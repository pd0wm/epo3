configuration timer_counter_timer_counter_arch_cfg of timer_counter is
   for timer_counter_arch
   end for;
end timer_counter_timer_counter_arch_cfg;


