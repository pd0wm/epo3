configuration score_tb_behaviour_cfg of score_tb is
   for behaviour
   end for;
end score_tb_behaviour_cfg;


