configuration debounce_testb_behaviour_cfg of debounce_testb is
   for behaviour
      for all: debounce use configuration work.debounce_behaviour_cfg;
      end for;
   end for;
end debounce_testb_behaviour_cfg;


