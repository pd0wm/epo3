configuration log_extracted_cfg of log is
   for extracted
   end for;
end log_extracted_cfg;


