configuration cs_shift_comb_cs_shift_comb_behav_cfg of cs_shift_comb is
   for cs_shift_comb_behav
   end for;
end cs_shift_comb_cs_shift_comb_behav_cfg;


