configuration vga_counter_8bitset_vga_counter_8bitset_behav_cfg of vga_counter_8bitset is
   for vga_counter_8bitset_behav
   end for;
end vga_counter_8bitset_vga_counter_8bitset_behav_cfg;


