configuration mux5_mux5_behav_cfg of mux5 is
   for mux5_behav
   end for;
end mux5_mux5_behav_cfg;


