configuration draw_score_behaviour_cfg of draw_score is
   for behaviour
   end for;
end draw_score_behaviour_cfg;


