configuration demux4_inv_demux4_inv_behav_cfg of demux4_inv is
   for demux4_inv_behav
   end for;
end demux4_inv_demux4_inv_behav_cfg;


