configuration debounce_tb_behaviour_cfg of debounce_tb is
   for behaviour
      for all: debounce use configuration work.debounce_behaviour_cfg;
      end for;
   end for;
end debounce_tb_behaviour_cfg;


