configuration vga_counter_3bit_vga_counter_3bit_behav_cfg of vga_counter_3bit is
   for vga_counter_3bit_behav
   end for;
end vga_counter_3bit_vga_counter_3bit_behav_cfg;


