configuration score_syn_tb_behaviour_cfg of score_tb is
   for behaviour
      for all: score use configuration work.score_synthesised_cfg;
      end for;
   end for;
end score_syn_tb_behaviour_cfg;


