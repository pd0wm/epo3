configuration controller_tb_controller_tb_arch_cfg of controller_tb is
   for controller_tb_arch
      for all: controller use configuration work.controller_controller_arch_cfg;
      end for;
   end for;
end controller_tb_controller_tb_arch_cfg;


