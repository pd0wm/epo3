configuration cs_7bc_cs_7bc_behav_cfg of cs_7bc is
   for cs_7bc_behav
   end for;
end cs_7bc_cs_7bc_behav_cfg;


