library IEEE;
use IEEE.std_logic_1164.ALL;

entity log_score_tb is
end log_score_tb;


