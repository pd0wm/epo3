library ieee;
use ieee.std_logic_1164.all;

package mem_params is
	constant mem_len : integer := 2**4;
	constant mem_addr_len : integer := 4;
	constant mem_subaddr_len : integer := 2;
end mem_params;

package body mem_params is
end mem_params;