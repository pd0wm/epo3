configuration rom_extracted_cfg of rom is
   for extracted
   end for;
end rom_extracted_cfg;


