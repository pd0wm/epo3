library IEEE;
use IEEE.std_logic_1164.ALL;

entity checkmask_tb is
end checkmask_tb;
