configuration cs_tri8_cs_tri8_behav_cfg of cs_tri8 is
   for cs_tri8_behav
   end for;
end cs_tri8_cs_tri8_behav_cfg;


