configuration vga_tb_vga_tb_arch_cfg2 of vga_tb is
   for vga_tb_arch
      for all: vga use configuration work.vga_extracted_cfg;
      end for;
   end for;
end vga_tb_vga_tb_arch_cfg2;


