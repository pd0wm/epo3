configuration vga_counter_2bit_vga_counter_2bit_behav_cfg of vga_counter_2bit is
   for vga_counter_2bit_behav
   end for;
end vga_counter_2bit_vga_counter_2bit_behav_cfg;


