configuration clearandshift_synthesised_cfg of clearandshift is
   for synthesised
   end for;
end clearandshift_synthesised_cfg;


