configuration vga_field_check_vga_field_check_arch_cfg of vga_field_check is
   for vga_field_check_arch
   end for;
end vga_field_check_vga_field_check_arch_cfg;


