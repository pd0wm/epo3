configuration controller_move_controller_move_arch_cfg of controller_move is
   for controller_move_arch
   end for;
end controller_move_controller_move_arch_cfg;


