configuration npg_mux2_1_behaviour_cfg of npg_mux2_1 is
   for behaviour
   end for;
end npg_mux2_1_behaviour_cfg;


