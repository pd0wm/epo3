configuration checkmask_tb_behaviour_syn_cfg of checkmask_tb is
   for checkmask_tb_behaviour
      for all: checkmask use configuration work.checkmask_synthesised_cfg;
      end for;
   end for;
end checkmask_tb_behaviour_syn_cfg;


