configuration tri_buff_extracted_cfg of tri_buff is
   for extracted
   end for;
end tri_buff_extracted_cfg;


