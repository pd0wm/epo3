configuration score_extr_tb_behaviour_cfg of score_tb is
   for behaviour
      for all: score use configuration work.score_extracted_cfg;
      end for;
   end for;
end score_extr_tb_behaviour_cfg;


