configuration vga_counter_8bit_vga_counter_8bit_behav_cfg of vga_counter_8bit is
   for vga_counter_8bit_behav
   end for;
end vga_counter_8bit_vga_counter_8bit_behav_cfg;


