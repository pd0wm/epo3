configuration piece_lut_behaviour_cfg of piece_lut is
   for piece_lut_behaviour
   end for;
end piece_lut_behaviour_cfg;


