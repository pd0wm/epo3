library IEEE;
use IEEE.std_logic_1164.ALL;

entity depiece_simple is
end depiece_simple;


