library IEEE;
use IEEE.std_logic_1164.ALL;

entity draw_score_tb is
end draw_score_tb;


