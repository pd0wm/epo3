configuration npg_tb_behaviour_cfg of npg_tb is
   for behaviour
      for all: npg use configuration work.npg_structural_cfg;
      end for;
   end for;
end npg_tb_behaviour_cfg;


