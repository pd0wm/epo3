configuration rom_mux4_behaviour_cfg of rom_mux4 is
   for rom_mux4_behaviour
   end for;
end rom_mux4_behaviour_cfg;


